/*
* Andrew Plaza
* Dr. Bishop
* VeriLog Assignment 3: Algorithmic Logic Unit
*/

`include "mux.v"

module alu;

endmodule
